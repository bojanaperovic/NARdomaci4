
module ram();

parameter size = 4096; // velicina rama u bitovima

reg [31:0] ram [0:size-1]; 

endmodule
